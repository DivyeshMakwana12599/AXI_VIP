//class ei_axi4_coverage_c 
  
//endclass : ei_axi4_coverage_c 
