hello

ddghad
dadadj
adsddd

