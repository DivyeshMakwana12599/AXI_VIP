//including all testcases files

`include "../test/ei_axi4_base_test.sv"
`include "../test/ei_axi4_read_test.sv"
`include "../test/ei_axi4_write_test.sv"
`include "../test/ei_axi4_sanity_test.sv"
`include "../test/ei_axi4_random_test.sv"
`include "../test/ei_axi4_seq_wr_rd_test.sv"
