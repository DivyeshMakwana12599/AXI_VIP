hello

ddghad
dadadj

