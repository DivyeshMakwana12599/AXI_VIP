`include "ei_axi4_macros.sv"
`include "ei_axi4_interface.sv"
`include "ei_axi4_assertion.sv"
`include "ei_axi4_coverage.sv"
`include "ei_axi4_checker.sv"
`include "ei_axi4_test_config.sv"
`include "ei_axi4_test.sv"
`include "ei_axi4_env_config.sv"
`include "ei_axi4_environment.sv"
`include "ei_axi4_transaction.sv"
`include "ei_axi4_reference_model.sv"
`include "ei_axi4_scoreboard.sv"
`include "ei_axi4_master_agent.sv"
`include "ei_axi4_slave_agent.sv"
`include "ei_axi4_master_generator.sv"
`include "ei_axi4_master_driver.sv"
`include "ei_axi4_master_transmit_monitor.sv"
`include "ei_axi4_slave_driver.sv"
`include "ei_axi4_slave_receive_monitor.sv"