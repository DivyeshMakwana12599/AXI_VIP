//including all testcases files

`include "../test/ei_axi4_base_test.sv"
// `include "../test/ei_axi4_read_test.sv"
// `include "../test/ei_axi4_write_test.sv"
`include "../test/ei_axi4_sanity_test.sv"
// `include "../test/ei_axi4_random_test.sv"
// `include "../test/ei_axi4_seq_wr_rd_test.sv"
// `include "../test/ei_axi4_4kb_boundary_test.sv"
// `include "../test/ei_axi4_parallel_wr_rd_test.sv"
// `include "../test/ei_axi4_error_wrap_unaligned_test.sv"
// `include "../test/ei_axi4_error_fixed_len_test.sv"
// `include "../test/ei_axi4_error_wrap_len_test.sv"
// `include "../test/ei_axi4_error_early_termination_test.sv"
