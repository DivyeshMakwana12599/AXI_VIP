`include "../src/ei_axi4_macros.sv"

`include "../src/ei_axi4_helper_functions.sv"

`include "../src/ei_axi4_transaction.sv"

`include "../src/ei_axi4_assertion.sv"

`include "../src/ei_axi4_coverage.sv"

`include "../src/ei_axi4_interface.sv"


`include "../src/ei_axi4_checker_cfg.sv"
`include "../src/ei_axi4_checker_db.sv"
`include "../src/ei_axi4_checker.sv"

`include "../test/ei_axi4_test_config.sv"
`include "../env/ei_axi4_env_config.sv"

`include "../src/ei_axi4_master_generator.sv"
`include "../src/ei_axi4_master_driver.sv"
`include "../src/ei_axi4_master_monitor.sv"
`include "../src/ei_axi4_master_agent.sv"

`include "../src/ei_axi4_slave_driver.sv"
`include "../src/ei_axi4_slave_monitor.sv"
`include "../src/ei_axi4_slave_agent.sv"

`include "../src/ei_axi4_reference_model.sv"
`include "../src/ei_axi4_scoreboard.sv"

`include "../env/ei_axi4_environment.sv"

`include "../test/ei_axi4_test.sv"
